module tt_um_priority_encoder (
    input  [7:0] A,      // Upper 8 bits
    input  [7:0] B,      // Lower 8 bits
    output reg [7:0] C   // Output position of the first '1'
);
    wire [15:0] In;      // Concatenated input

    assign In = {A, B};  // In[15:0] = {A[7:0], B[7:0]}

    always @(*) begin
        casez (In)  
            16'b1???????????????: C = 8'd15;
            16'b01??????????????: C = 8'd14;
            16'b001?????????????: C = 8'd13;
            16'b0001????????????: C = 8'd12;
            16'b00001???????????: C = 8'd11;
            16'b000001??????????: C = 8'd10;
            16'b0000001?????????: C = 8'd9;
            16'b00000001????????: C = 8'd8;
            16'b000000001???????: C = 8'd7;
            16'b0000000001??????: C = 8'd6;
            16'b00000000001?????: C = 8'd5;
            16'b000000000001????: C = 8'd4;
            16'b0000000000001???: C = 8'd3;
            16'b00000000000001??: C = 8'd2;
            16'b000000000000001?: C = 8'd1;
            16'b0000000000000001: C = 8'd0;
            16'b0000000000000000: C = 8'b11110000; // Special case
            default: C = 8'b00000000;
        endcase
    end
endmodule